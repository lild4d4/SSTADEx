** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/SSTADEx/test/sstadex/xschem/ldo_sim_ihp.sch
**.subckt ldo_sim_ihp
I2 vs vss 40e-6
I1 vmid vss 20e-6
C8 vout_s1 vmid 3e-12 m=1
R1 vout vfb 100000 m=1
R2 vfb vss 300000 m=1
Cl vout vss 10e-9 m=1
R3 vout vss 18 m=1
XM1 vout_s1 vfb vs vs sg13_hv_nmos w=2.13u l=0.8u ng=1 m=1
XM2 net1 vn vs vs sg13_hv_nmos w=2.13u l=0.8u ng=1 m=1
XM3 vout_s1 net1 vdd vdd sg13_hv_pmos w=0.41u l=0.4u ng=1 m=1
XM4 net1 net1 vdd vdd sg13_hv_pmos w=0.41u l=0.4u ng=1 m=1
XM5 vmid vout_s1 vdd vdd sg13_hv_pmos w=0.41u l=0.4u ng=1 m=1
XM6 vout vmid vdd vdd sg13_hv_pmos w=2487u l=0.4u ng=1 m=1
**** begin user architecture code



.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOShv.lib mos_tt

Vref vn 0 1.35
Vdd vdd 0 3.3 ac 1
Vss vss 0 0

.control
pre_osdi /opt/pdks/ihp-sg13g2/libs.tech/ngspice/openvaf/psp103_nqs.osdi
ac dec 10 1 100G
let gm_diff = @n.xm1.nsg13_hv_nmos[gm]
let gds_diff = @n.xm1.nsg13_hv_nmos[gds]
let gm_al = @n.xm3.nsg13_hv_pmos[gm]
let gds_al = @n.xm3.nsg13_hv_pmos[gds]
wrdata temp.csv vdb(vout) phase(vout) gm_diff gds_diff gm_al gds_al v(vout)
.endc



**** end user architecture code
**.ends
.end