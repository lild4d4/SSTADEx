** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/SSTADEx/test/Tesis_notebooks/xschem/ota_2stage_tb.sch
**.subckt ota_2stage_tb
XM1 vout_s1 vn vs vs sg13_hv_nmos L=3.1999999999999997u W=309.4677996593u ng=1 m=1 
XM2 net2 net1 vs vs sg13_hv_nmos L=3.1999999999999997u W=309.4677996593u ng=1 m=1 
XM3 vout_s1 net2 vdd vdd sg13_hv_pmos L=6.3999999999999995u W=177.8724061624u ng=1 m=1 
XM4 net2 net2 vdd vdd sg13_hv_pmos L=6.3999999999999995u W=177.8724061624u ng=1 m=1 
XM5 vout vout_s1 vdd vdd sg13_hv_pmos L=3.1999999999999997u W=170.474533378u ng=1 m=1 
R1 vfb vout 10000000000 m=1
C2 vfb vss 10 m=1
R2 vfb vss -42857142857 m=1
V1 net1 vfb dc 0 ac 1
C3 vout vss 2.026e-11 m=1
XM6 vss net3 vs vss sg13_hv_nmos L=6.3999999999999995u W=54.14271527541397u ng=1 m=1 
XM7 vss net3 net3 vss sg13_hv_nmos L=6.3999999999999995u W=54.14271527541397u ng=1 m=1 
I2 vdd net3 4e-05 
XM8 vss net3 vout vss sg13_hv_nmos L=6.3999999999999995u W=54.14271527541397u ng=1 m=1 
Cc vout_s1 net4 1e-10 m=1 
Rc vout net4 10000.0 m=1 
**** begin user architecture code



.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOShv.lib mos_tt

Vref vn 0 0.9
Vdd vdd 0 1.8
Vss vss 0 0

.control
pre_osdi /opt/pdks/ihp-sg13g2/libs.tech/ngspice/openvaf/psp103_nqs.osdi
ac dec 10 1 1G
wrdata temp.csv vdb(vout) phase(vout)
.endc