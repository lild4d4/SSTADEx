** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/SSTADEx/test/sstadex/xschem/stage2_OTA_tb_ihp.sch
**.subckt stage2_OTA_tb_ihp
I2 vs vss 40e-6
I1 vout vss 20e-6
C1 vout vss 1e-12 m=1
XM1 vout_s1 vn vs vs sg13_hv_nmos w=219.27u l=0.8u ng=1 m=1
XM2 net2 net1 vs vs sg13_hv_nmos w=219.27u l=0.8u ng=1 m=1
XM3 vout_s1 net2 vdd vdd sg13_hv_pmos w=10.48u l=0.4u ng=1 m=1
XM4 net2 net2 vdd vdd sg13_hv_pmos w=10.48u l=0.4u ng=1 m=1
XM5 vout vout_s1 vdd vdd sg13_hv_pmos w=31.32u l=0.8u ng=1 m=1
R1 vfb vout 100000000 m=1
C2 vfb vss 10 m=1
R2 vfb vss 450000000 m=1
V1 net1 vfb dc 0 ac 1
**** begin user architecture code



.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOShv.lib mos_tt

Vref vn 0 1.35
Vdd vdd 0 3.3
Vss vss 0 0

.param vcc=3.3

.control
pre_osdi /opt/pdks/ihp-sg13g2/libs.tech/ngspice/openvaf/psp103_nqs.osdi
ac dec 10 1 1G
let gm_diff = @n.xm1.nsg13_hv_nmos[gm]
let gds_diff = @n.xm1.nsg13_hv_nmos[gds]
let gm_al = @n.xm3.nsg13_hv_pmos[gm]
let gds_al = @n.xm3.nsg13_hv_pmos[gds]
wrdata temp.csv vdb(vout) phase(vout) gm_diff gds_diff gm_al gds_al v(vout)
.endc



**** end user architecture code
**.ends
.end