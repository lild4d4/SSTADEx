** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/SSTADEx/test/Tesis_notebooks/xschem/ldo_ol_cap.sch
**.subckt ldo_ol_cap
Gdif_m1_1 net1 vss net2 vss 0.0001414
Raload_m1_1 vss net3 6.5283e4 m=1
Gaload_m1_1 net3 vss net4 vss 1.47e-5
Gdif_m2_1 net4 net1 vss net1 6.97e-5
Ccpdif vss net1 9e-13 m=1
Raload_m2_1 net3 net4 3.328e6 m=1
Gaload_m2_1 net4 net3 vss net3 2.5e-4
Ccpaload_m1 net4 net3 5.74e-14 m=1
Ccpaload_m2 net3 vss 3.2e-12 m=1
R1 vout vfb 5000 m=1
R2 vfb vss 15000 m=1
Ro_pt vss vout 202 m=1
Gm_pt vout vss net4 vss 0.1860
Cgg_pt net4 vss 1.59e-12 m=1
Cgd_pt net4 vout 8.6e-15 m=1
R4 vpos vfb 10000000000 m=1
C2 vpos vss 10 m=1
V1 net2 vpos dc 0 ac 1
Cl vout vss 1e-12 m=1
R3 vout vss 18 m=1
Ca net4 vss 7.37e-10 m=1
Rdif_1 net1 vss 82143691 m=1
Rdif_2 net4 net1 82143691 m=1
**** begin user architecture code



.lib /opt/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt

Vss vss 0 0

.control
ac dec 10 1 10G
plot vdb(vout)
plot phase(vout)*180/PI
.endc



**** end user architecture code
**.ends
.end
