** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/SSTADEx/test/Tesis_notebooks/xschem/ota_1stage_tb.sch
**.subckt ota_1stage_tb
XM1 vs net1 vout vs sg13_hv_nmos w=100.4u l=0.45u ng=1 m=1
XM2 vs vn net2 vs sg13_hv_nmos w=100.4u l=0.45u ng=1 m=1
XM3 vout net2 vdd vdd sg13_hv_pmos w=10.48u l=0.4u ng=1 m=1
XM4 net2 net2 vdd vdd sg13_hv_pmos w=10.48u l=0.4u ng=1 m=1
R1 vfb vout 10000000000 m=1
C2 vfb vss 10 m=1
R2 vfb vss 90000000000 m=1
XM5 vss net3 vs vss sg13_hv_nmos w=34.32u l=0.45u ng=1 m=1
XM6 vss net3 net3 vss sg13_hv_nmos w=34.32u l=0.45u ng=1 m=1
I2 vdd net3 40e-6
V1 net1 vfb dc 0 ac 1
**** begin user architecture code



.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOShv.lib mos_tt

Vref vn 0 0.9
Vdd vdd 0 1.8
Vss vss 0 0

.control
ac dec 10 1 1G
plot vdb(vout)
plot phase(vout)
op
print vout vs vfb
.endc



**** end user architecture code
**.ends
.end
