** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/SSTADEx/test/Tesis_notebooks/xschem/mna_example.sch
**.subckt mna_example
R1 vout vss 1 m=1
G1 vout vss net2 net3 1e-6
C1 vout vss 1 m=1
I0 vdd vout 1m
C2 net1 vss 1 m=1
C3 net1 vout 1 m=1
V1 net1 vss 3
**.ends
.end
