* Lookup Table Generation *
.lib '/opt/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt'
VGS NG 0 DC=0
VBS NB 0 DC=0
VDS ND 0 DC=0
XM1 ND NG 0 NB sky130_fd_pr__nfet_01v8 L=0.6 W=20.0

.options TEMP = 27
.options TNOM = 27
.control
save i(vds)
dc VDS 0.0 3.3 0.01 VGS 0.0 3.3 0.01
let i_vds = abs(i(vds))
write /tmp/tmp23te_z82 all
.endc
.end