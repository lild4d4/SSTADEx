** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/SSTADEx/test/Tesis_notebooks/xschem/ota_2stage_v2.sch
**.subckt ota_2stage_v2
Ro_2stage vdd vout 100 m=1
Gm_2stage vout vdd vin vdd 1
V1 vdd vss 1
Cin_2stage vin vdd 1e-12 m=1
V2 vin vss 1
Gcs_2stage vout vss vss vss 1
Rcs_2stage vss vout 100 m=1
Cin_pt vout vss 1e-12 m=1
**.ends
.end