** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/SSTADEx/test/Tesis_notebooks/xschem/ldo_tb.sch
**.subckt ldo_tb
R1 vout vfb 22500 m=1
R2 vfb vss 67500 m=1
Cl vout vss 1e-12 m=1
XM1 vout_s1 vfb vs vs sg13_hv_nmos w=5.33u l=0.8u ng=1 m=1
XM2 net1 vn vs vs sg13_hv_nmos w=5.33u l=0.8u ng=1 m=1
XM3 vout_s1 net1 vdd_1 vdd_1 sg13_hv_pmos w=9.02u l=6.4u ng=1 m=1
XM4 net1 net1 vdd_1 vdd_1 sg13_hv_pmos w=9.02u l=6.4u ng=1 m=1
XM5 vmid vout_s1 vdd_1 vdd_1 sg13_hv_pmos w=8.8u l=3.2u ng=1 m=1
XM9 vout vmid vdd vdd sg13_hv_pmos w=2488u l=0.4u ng=1 m=1
R3 vout vss 18 m=1
XM6 vss net2 vs vss sg13_hv_nmos w=5.4u l=3.2u ng=1 m=1
XM7 vss net2 net2 vss sg13_hv_nmos w=5.4u l=3.2u ng=1 m=1
XM8 vss net2 vmid vss sg13_hv_nmos w=5.4u l=3.2u ng=1 m=1
I2 vdd_1 net2 40e-6
**** begin user architecture code



.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOShv.lib mos_tt

Vref vn 0 1.35
Vdd vdd 0 3.3 ac 1
Vdd_1 vdd_1 0 3.3
Vss vss 0 0

.control
pre_osdi /opt/pdks/ihp-sg13g2/libs.tech/ngspice/openvaf/psp103_nqs.osdi
ac dec 10 1 1G
wrdata temp.csv vdb(vout) phase(vout)
.endc



**** end user architecture code
**.ends
.end