* sch_path: /workspaces/usm-vlsi-tools/shared_xserver/SSTADEx/test/Tesis_notebooks/xschem/ota_tb_ihp_cc_full.sch
**.subckt ota_tb_ihp_cc_full
I2 vs vss 20e-6
XM1 vcp vp1 vs vs sg13_hv_nmos w=5.4u l=0.4u ng=1 m=1
XM2 net2 vn vs vs sg13_hv_nmos w=5.4u l=0.4u ng=1 m=1
XM3 vout vbias_dp vcp vcp sg13_hv_nmos w=5.8u l=0.8u ng=1 m=1
XM4 net1 vbias_dp net2 net2 sg13_hv_nmos w=5.8u l=0.8u ng=1 m=1
XM5 net3 net1 vdd vdd sg13_hv_pmos w=5.5u l=6.4u ng=1 m=1
XM6 vcp_cm net1 vdd vdd sg13_hv_pmos w=5.5u l=6.4u ng=1 m=1
R1 vfb vout 10000000000 m=1
C2 vfb vss 10 m=1
R2 vfb vss 38571428570 m=1
V1 vp1 vfb dc 0 ac 1
XM7 net1 vbias_cm net3 net3 sg13_hv_pmos w=5.2u l=0.8u ng=1 m=1
XM8 vout vbias_cm vcp_cm vcp_cm sg13_hv_pmos w=5.2u l=0.8u ng=1 m=1
**** begin user architecture code



.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOShv.lib mos_tt

Vref vn 0 1.35
Vdd vdd 0 3.3
Vbias_dp vbias_dp 0 2.2
Vbias_cm vbias_cm vdd -2.1
Vss vss 0 0

.control
pre_osdi /opt/pdks/ihp-sg13g2/libs.tech/ngspice/openvaf/psp103_nqs.osdi
ac dec 10 1 1G
*plot vdb(vout)
*plot phase(vout)*180/PI
*meas ac gain find vdb(vout) at=1
*let low_gain = gain-3
*meas ac fc WHEN vdb(vout)=low_gain
wrdata temp.csv vdb(vout) phase(vout)
.endc



**** end user architecture code
**.ends
.end