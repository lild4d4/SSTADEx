** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/AC3E-IHP_ALDO/xschem/ota/ota_tb_openloop.sch
**.subckt ota_tb_openloop
V1 vcm vss DC{vcm}
V2 vsen vcm sin(0 {vac} 1Meg) dc 0 ac 1
V4 vdd vss DC {vdd}
V5 vss GND DC{vss}
I0 vss net1 DC{iref}
R1 net3 vcm 500 m=1
C2 vin vsen 1 m=1
R2 vout net2 5k m=1
C3 vout vss 10p m=1
R3 vin net2 1G m=1
x1 vin vcm net1 vdd vss vout ota
**** begin user architecture code


.param iref = 5u
.param vdd  = 1.8
.param vss  = 0.0
.param vcm  = 0.9
.param vac  = 60m

* OP Parameters & Singals to save


*Simulation

.control
reset
*pre_osdi /opt/pdks/ihp-sg13g2/libs.tech/ngspice/openvaf/psp103_nqs.osdi
set color0 = white
ac dec 100 1 10G
remzerovec
write ota_tb_openloop_ac.raw
setplot ac1
meas ac GBW when vdb(vout)=0
meas ac DCG find vdb(vout) at=1
meas ac PM find vp(vout) when vdb(vout)=0
print PM*180/PI
meas ac GM find vdb(vout) when vp(vout)=0
wrdata ota_tb_openloop_ac.csv vdb(vout) {vp(vout)*180/PI}

.endc

*.control
*tran 1e-6 1e-3
*write test_tran.raw
*noise V(vout) V2 dec 10 10 100e3
*print inoise_total onoise_total
*.endc

*.control
*alter V2 ac 0
*alter v4 ac 1
*tran 1e-6 1e-3
*write test_tran.raw
*noise V(vout) V4 dec 10 10 100e3
*print inoise_total onoise_total
*.endc

.end




.param corner=0

.if (corner==0)
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ
.endif

**** end user architecture code
**.ends

* expanding   symbol:  /workspaces/usm-vlsi-tools/shared_xserver/AC3E-IHP_ALDO/xschem/ota/ota.sym # of pins=6
** sym_path: /workspaces/usm-vlsi-tools/shared_xserver/AC3E-IHP_ALDO/xschem/ota/ota.sym
** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/AC3E-IHP_ALDO/xschem/ota/ota.sch
.subckt ota vin_n vin_p iref vdd vss vout
*.ipin iref
*.ipin vin_n
*.ipin vin_p
*.iopin vdd
*.iopin vss
*.opin vout
XM1 net1 vin_n net2 vss sg13_lv_nmos w=15u l=2u ng=1 m=1
XM2 net3 vin_p net2 vss sg13_lv_nmos w=15u l=2u ng=1 m=1
XM3 net3 net1 vdd vdd sg13_lv_pmos w=2u l=1u ng=1 m=1
XM4 net1 net1 vdd vdd sg13_lv_pmos w=2u l=1u ng=1 m=1
XM5 net2 iref vss vss sg13_lv_nmos w=6u l=2u ng=1 m=1
XM8 iref iref vss vss sg13_lv_nmos w=6u l=2u ng=1 m=1
XM6 vout net3 vdd vdd sg13_lv_pmos w=20u l=0.5u ng=1 m=1
XM7 vout iref vss vss sg13_lv_nmos w=24u l=2u ng=1 m=1
XR2 net3 net4 rhigh w=0.5e-6 l=10e-6 m=1 b=0
XC2 net4 vout cap_cmim w=45.0e-6 l=45.0e-6 m=1
.ends

.GLOBAL GND
.end
