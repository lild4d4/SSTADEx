** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/SSTADEx/test/Tesis_notebooks/untitled.sch
**.subckt untitled
R3 vpos vfb 100000000 m=1
C1 vpos vss 10 m=1
Ro_pt vss vout 1314 m=1
Gm_pt vout vss net1 vss 0.225
R1 vout vfb 328 m=1
R2 vfb vss 984 m=1
Gma net1 vss vss vol 0.01
Ra vss net1 10000000 m=1
Rl vout vss 12 m=1
Cgg_pt net1 vss 1.86e-11 m=1
Ca net1 vss 1e-17 m=1
Cl vout vss 1e-12 m=1
V3 vol vpos dc 0 ac 1
Cgg_pt1 net1 vout 1.86e-14 m=1
**** begin user architecture code



Vss vss 0 0

.control

ac dec 10 1 1G
plot vdb(vout)
plot phase(vout)*180/PI


.endc



**** end user architecture code
**.ends
.end
