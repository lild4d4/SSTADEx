** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/SSTADEx/test/Tesis_notebooks/xschem/ldo_ol_sim_ihp_cc.sch
**.subckt ldo_ol_sim_ihp_cc
R1 vout vfb 100000 m=1
R2 vfb vss 300000 m=1
Cl vout vss 1e-12 m=1
R3 vout vss 18 m=1
XM6 vmid net2 vdd vdd sg13_hv_pmos w=10.97u l=6.4u ng=1 m=1
I2 vs vss 40e-6
XM1 vcp vn vs vs sg13_hv_nmos w=5.87u l=6.4u ng=1 m=1
XM2 net3 net1 vs vs sg13_hv_nmos w=5.87u l=6.4u ng=1 m=1
XM3 vmid vbias vcp vcp sg13_hv_nmos w=6.42u l=0.8u ng=1 m=1
XM4 net2 vbias net3 net3 sg13_hv_nmos w=6.42u l=0.8u ng=1 m=1
XM5 net2 net2 vdd vdd sg13_hv_pmos w=10.97u l=6.4u ng=1 m=1
XM7 vout vmid vdd vdd sg13_hv_pmos w=2487u l=0.4u ng=1 m=1
R4 vpos vfb 100000000 m=1
C2 vpos vss 10 m=1
V1 net1 vpos dc 0 ac 1
Cl1 vmid vout 3e-12 m=1
**** begin user architecture code



.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOShv.lib mos_tt

Vref vn 0 1.35
Vdd vdd 0 3.3
Vss vss 0 0
Vbias vbias 0 2.2

.control
ac dec 10 1 100G
plot vdb(vout)
plot phase(vout)*180/PI
op
print vout vmid vcp vfb vs
.endc



**** end user architecture code
**.ends
.end
